module deathROM(input [7:0] addr,
                output [15:0] data);

    parameter ADDR_WIDTH = 8;
    parameter DATA_WIDTH = 16;
	
    parameter [0:2**ADDR_WIDTH - 1][DATA_WIDTH-1:0] ROM = {
            //code x00 - pacman closed
        16'b0000000000000000, // 0
        16'b0000011111000000, // 1
        16'b0001111111110000, // 2
        16'b0011111111111000, // 3
        16'b0011111111111000, // 4
        16'b0111111111111100, // 5
        16'b0111111111111100, // 6
        16'b0111111111111100, // 7
        16'b0111111111111100, // 8
        16'b0111111111111100, // 9
        16'b0011111111111000, // 10
        16'b0011111111111000, // 11
        16'b0001111111110000, // 12
        16'b0000011111000000, // 13
        16'b0000000000000000, // 14
        16'b0000000000000000, // 15
            //code x01 - death one 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0110000000001100,
        16'b0111000000011100,
        16'b0111100000111100,
        16'b0111110001111100,
        16'b0111111011111100,
        16'b0011111111111000,
        16'b0011111111111000,
        16'b0001111111110000,
        16'b0000011111000000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x02 - death two 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0100000000000100,
        16'b1111000000011110,
        16'b1111100000111110,
        16'b1111111011111110,
        16'b0111111111111100,
        16'b0111111111111100,
        16'b0011111111111000,
        16'b0000111011100000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x03 - death three 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b1110000000001110,
        16'b1111110001111110,
        16'b1111111111111110,
        16'b0111111111111100,
        16'b0011111111111000,
        16'b0000111011100000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x04 - death four 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b1111000000011110,
        16'b1111111111111110,
        16'b1111111111111110,
        16'b0111111111111100,
        16'b0001111011110000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x05 - death five
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000111111100000,
        16'b1111111111111110,
        16'b1111111111111110,
        16'b0111111111111100,
        16'b0001111011110000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x06 - death six 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000001110000000,
        16'b0000111111100000,
        16'b0111111111111100,
        16'b1111111111111110,
        16'b0111111011111100,
        16'b0001110001110000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x07 - death seven 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000100000000,
        16'b0000001110000000,
        16'b0000111111100000,
        16'b0001111111110000,
        16'b0111111111111100,
        16'b0111111011111100,
        16'b0011110001111000,
        16'b0000000000000000,
            //code x08 - death eight 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000100000000,
        16'b0000001110000000,
        16'b0000011111000000,
        16'b0000011111000000,
        16'b0000111111100000,
        16'b0001111111110000,
        16'b0000111011100000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x09 - death nine 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000100000000,
        16'b0000000100000000,
        16'b0000001110000000,
        16'b0000001110000000,
        16'b0000001110000000,
        16'b0000011111000000,
        16'b0000001010000000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x0A - death ten 
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000100000000,
        16'b0000000100000000,
        16'b0000000100000000,
        16'b0000000100000000,
        16'b0000000100000000,
        16'b0000000100000000,
        16'b0000000000000000,
        16'b0000000000000000,
            //code x0B - death eleven
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000010001000000,
        16'b0001001010000000,
        16'b0000100000010000,
        16'b0000000000100000,
        16'b0011000000000000,
        16'b0000000000011000,
        16'b0000100000000000,
        16'b0001000000100000,
        16'b0000001010010000,
        16'b0000010001000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000
    };
    assign data = ROM[addr]; 
endmodule 