//         
//			// code x41
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00010000, // 2    *
//        8'b00111000, // 3   ***
//        8'b01101100, // 4  ** **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11111110, // 7 *******
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b11000110, // b **   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x42
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111100, // 2 ******
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01111100, // 6  *****
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11111100, // b ******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x43
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b01100110, // 3  **  **
//        8'b11000010, // 4 **    *
//        8'b11000000, // 5 **
//        8'b11000000, // 6 **
//        8'b11000000, // 7 **
//        8'b11000000, // 8 **
//        8'b11000010, // 9 **    *
//        8'b01100110, // a  **  **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x44
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111000, // 2 *****
//        8'b01101100, // 3  ** **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01100110, // 6  **  **
//        8'b01100110, // 7  **  **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01101100, // a  ** **
//        8'b11111000, // b *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x45
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111110, // 2 *******
//        8'b01100110, // 3  **  **
//        8'b01100010, // 4  **   *
//        8'b01101000, // 5  ** *
//        8'b01111000, // 6  ****
//        8'b01101000, // 7  ** *
//        8'b01100000, // 8  **
//        8'b01100010, // 9  **   *
//        8'b01100110, // a  **  **
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x46
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111110, // 2 *******
//        8'b01100110, // 3  **  **
//        8'b01100010, // 4  **   *
//        8'b01101000, // 5  ** *
//        8'b01111000, // 6  ****
//        8'b01101000, // 7  ** *
//        8'b01100000, // 8  **
//        8'b01100000, // 9  **
//        8'b01100000, // a  **
//        8'b11110000, // b ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x47
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b01100110, // 3  **  **
//        8'b11000010, // 4 **    *
//        8'b11000000, // 5 **
//        8'b11000000, // 6 **
//        8'b11011110, // 7 ** ****
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b01100110, // a  **  **
//        8'b00111010, // b   *** *
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x48
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000110, // 2 **   **
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11111110, // 6 *******
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b11000110, // b **   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x49
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00111100, // 2   ****
//        8'b00011000, // 3    **
//        8'b00011000, // 4    **
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4a
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b00011110, // 2    ****
//        8'b00001100, // 3     **
//        8'b00001100, // 4     **
//        8'b00001100, // 5     **
//        8'b00001100, // 6     **
//        8'b00001100, // 7     **
//        8'b11001100, // 8 **  **
//        8'b11001100, // 9 **  **
//        8'b11001100, // a **  **
//        8'b01111000, // b  ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4b
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11100110, // 2 ***  **
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01101100, // 5  ** **
//        8'b01111000, // 6  ****
//        8'b01111000, // 7  ****
//        8'b01101100, // 8  ** **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11100110, // b ***  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4c
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11110000, // 2 ****
//        8'b01100000, // 3  **
//        8'b01100000, // 4  **
//        8'b01100000, // 5  **
//        8'b01100000, // 6  **
//        8'b01100000, // 7  **
//        8'b01100000, // 8  **
//        8'b01100010, // 9  **   *
//        8'b01100110, // a  **  **
//        8'b11111110, // b *******
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4d
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11100111, // 3 ***  ***
//        8'b11111111, // 4 ********
//        8'b11111111, // 5 ********
//        8'b11011011, // 6 ** ** **
//        8'b11000011, // 7 **    **
//        8'b11000011, // 8 **    **
//        8'b11000011, // 9 **    **
//        8'b11000011, // a **    **
//        8'b11000011, // b **    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4e
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000110, // 2 **   **
//        8'b11100110, // 3 ***  **
//        8'b11110110, // 4 **** **
//        8'b11111110, // 5 *******
//        8'b11011110, // 6 ** ****
//        8'b11001110, // 7 **  ***
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b11000110, // b **   **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x4f
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x50
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111100, // 2 ******
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01111100, // 6  *****
//        8'b01100000, // 7  **
//        8'b01100000, // 8  **
//        8'b01100000, // 9  **
//        8'b01100000, // a  **
//        8'b11110000, // b ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x510
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11010110, // 9 ** * **
//        8'b11011110, // a ** ****
//        8'b01111100, // b  *****
//        8'b00001100, // c     **
//        8'b00001110, // d     ***
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x52
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111100, // 2 ******
//        8'b01100110, // 3  **  **
//        8'b01100110, // 4  **  **
//        8'b01100110, // 5  **  **
//        8'b01111100, // 6  *****
//        8'b01101100, // 7  ** **
//        8'b01100110, // 8  **  **
//        8'b01100110, // 9  **  **
//        8'b01100110, // a  **  **
//        8'b11100110, // b ***  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x53
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b01111100, // 2  *****
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b01100000, // 5  **
//        8'b00111000, // 6   ***
//        8'b00001100, // 7     **
//        8'b00000110, // 8      **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x54
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111111, // 2 ********
//        8'b11011011, // 3 ** ** **
//        8'b10011001, // 4 *  **  *
//        8'b00011000, // 5    **
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x55
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000110, // 2 **   **
//        8'b11000110, // 3 **   **
//        8'b11000110, // 4 **   **
//        8'b11000110, // 5 **   **
//        8'b11000110, // 6 **   **
//        8'b11000110, // 7 **   **
//        8'b11000110, // 8 **   **
//        8'b11000110, // 9 **   **
//        8'b11000110, // a **   **
//        8'b01111100, // b  *****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x56
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b11000011, // 4 **    **
//        8'b11000011, // 5 **    **
//        8'b11000011, // 6 **    **
//        8'b11000011, // 7 **    **
//        8'b11000011, // 8 **    **
//        8'b01100110, // 9  **  **
//        8'b00111100, // a   ****
//        8'b00011000, // b    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x57
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b11000011, // 4 **    **
//        8'b11000011, // 5 **    **
//        8'b11000011, // 6 **    **
//        8'b11011011, // 7 ** ** **
//        8'b11011011, // 8 ** ** **
//        8'b11111111, // 9 ********
//        8'b01100110, // a  **  **
//        8'b01100110, // b  **  **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//        
//         // code x58
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b01100110, // 4  **  **
//        8'b00111100, // 5   ****
//        8'b00011000, // 6    **
//        8'b00011000, // 7    **
//        8'b00111100, // 8   ****
//        8'b01100110, // 9  **  **
//        8'b11000011, // a **    **
//        8'b11000011, // b **    **
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x59
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11000011, // 2 **    **
//        8'b11000011, // 3 **    **
//        8'b11000011, // 4 **    **
//        8'b01100110, // 5  **  **
//        8'b00111100, // 6   ****
//        8'b00011000, // 7    **
//        8'b00011000, // 8    **
//        8'b00011000, // 9    **
//        8'b00011000, // a    **
//        8'b00111100, // b   ****
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f
//         // code x5aa
//        8'b00000000, // 0
//        8'b00000000, // 1
//        8'b11111111, // 2 ********
//        8'b11000011, // 3 **    **
//        8'b10000110, // 4 *    **
//        8'b00001100, // 5     **
//        8'b00011000, // 6    **
//        8'b00110000, // 7   **
//        8'b01100000, // 8  **
//        8'b11000001, // 9 **     *
//        8'b11000011, // a **    **
//        8'b11111111, // b ********
//        8'b00000000, // c
//        8'b00000000, // d
//        8'b00000000, // e
//        8'b00000000, // f