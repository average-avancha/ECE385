module ghostROM (input [7:0] addr,
                 output [63:0] data);
    parameter ADDR_WIDTH = 8;
    parameter DATA_WIDTH = 64;
	 
    parameter [0:2**ADDR_WIDTH - 1][DATA_WIDTH-1:0] ROM = {
		//x00 ghost open scared
		64'h0000000000000000,
		64'h0000001111000000,
		64'h0000111111110000,
		64'h0001111111111000,
		64'h0011111111111100,
		64'h0011111111111100,
		64'h0011133113311100,
		64'h0111133113311110,
		64'h0111111111111110,
		64'h0111111111111110,
		64'h0113311331133110,
		64'h0131133113311310,
		64'h0111111111111110,
		64'h0110111001110110,
		64'h0100011001100010,
		64'h0000000000000000,
		//x01 ghost close scared
		64'h0000000000000000,
		64'h0000001111000000,
		64'h0000111111110000,
		64'h0001111111111000,
		64'h0011111111111100,
		64'h0011111111111100,
		64'h0011133113311100,
		64'h0111133113311110,
		64'h0111111111111110,
		64'h0111111111111110,
		64'h0113311331133110,
		64'h0131133113311310,
		64'h0111111111111110,
		64'h0111101111011110,
		64'h0011000110001100,
		64'h0000000000000000,
		//x02 ghost open up
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000112222110000,
		64'h000a11a22a11a000,
		64'h002aaaa22aaaa200,
		64'h002aaaa22aaaa200,
		64'h0022aa2222aa2200,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0220222002220220,
		64'h0200022002200020,
		64'h0000000000000000,
		//x03 ghost close up
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000112222110000,
		64'h000a11a22a11a000,
		64'h002aaaa22aaaa200,
		64'h002aaaa22aaaa200,
		64'h0022aa2222aa2200,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222202222022220,
		64'h0022000220002200,
		64'h0000000000000000,
		//x04 ghost open left
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000222222220000,
		64'h0002222222222000,
		64'h002aa2222aa22200,
		64'h00aaaa22aaaa2200,
		64'h0011aa2211aa2200,
		64'h0211aa2211aa2220,
		64'h022aa2222aa22220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0220222002220220,
		64'h0200022002200020,
		64'h0000000000000000,
		//x05 ghost close left
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000222222220000,
		64'h0002222222222000,
		64'h002aa2222aa22200,
		64'h00aaaa22aaaa2200,
		64'h0011aa2211aa2200,
		64'h0211aa2211aa2220,
		64'h022aa2222aa22220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222202222022220,
		64'h0022000220002200,
		64'h0000000000000000,
		//x06 ghost open down
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000222222220000,
		64'h0002222222222000,
		64'h0022222222222200,
		64'h0022aa2222aa2200,
		64'h002aaaa22aaaa200,
		64'h022aaaa22aaaa220,
		64'h022a11a22a11a220,
		64'h0222112222112220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0220222002220220,
		64'h0200022002200020,
		64'h0000000000000000,
		//x07 ghost close down
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000222222220000,
		64'h0002222222222000,
		64'h0022222222222200,
		64'h0022aa2222aa2200,
		64'h002aaaa22aaaa200,
		64'h022aaaa22aaaa220,
		64'h022a11a22a11a220,
		64'h0222112222112220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222202222022220,
		64'h0022000220002200,
		64'h0000000000000000,
		//x08 ghost open right
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000222222220000,
		64'h0002222222222000,
		64'h00222aa2222aa200,
		64'h0022aaaa22aaaa00,
		64'h0022aa1122aa1100,
		64'h0222aa1122aa1120,
		64'h02222aa2222aa220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0220222002220220,
		64'h0200022002200020,
		64'h0000000000000000,
		//x09 ghost close right
		64'h0000000000000000,
		64'h0000002222000000,
		64'h0000222222220000,
		64'h0002222222222000,
		64'h00222AA2222AA200,
		64'h0022AAAA22AAAA00,
		64'h0022AA1122AA1100,
		64'h0222AA1122AA1120,
		64'h02222AA2222AA220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222222222222220,
		64'h0222202222022220,
		64'h0022000220002200,
		64'h0000000000000000
	 };
    assign data = ROM[addr]; 
endmodule 