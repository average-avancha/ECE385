//module pacman_spriteFSM(input        Clk, frame_clk_rising_edge,
//                        input        Reset,
//                        input        increment_score_powdot,
//                        output [4:0] timer_powered_up,
//                        output       pac_powered_up);
//
//endmodule 
