module mapROM_parallel(input  [8:0] addr, 
							  output [511:0] data [0:15]);
	 parameter ADDR_WIDTH = 9;
    parameter DATA_WIDTH = 512;
	 
	 parameter [0:2**ADDR_WIDTH - 1][DATA_WIDTH-1:0] ROM = {
		512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
		512'b11010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011,
		512'b10010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001,
		512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000011111111111111111111111111111100000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000011111111111111111111111111111100000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000111111111111111111111111110000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000001111111111111111111111111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000011000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000011000000000000000000000000111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000001111111111111111111111111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000111100000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000011000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111110000000000000000000111100000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000111100000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000001100000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000111100000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000111100000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000111100000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000111100000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000111100000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000111100000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000111100000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000111100000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000111100000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000111100000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000000111111111100000000000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000000001111111111111100000000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000011111111111111111000000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000000111111111111111111000000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000001111111111111111111100000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000001111111111111111111100000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000011111111111111111111110000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000011111111111111111111110000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000001111111111111111111111110000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111100000000000000000000000000011111111111111111111110000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111110000000000000000011111111111111111111111110000000000000000000000000001111111111110000000000000000000111100000000000000000001111111111111100000000000000000000000000011111111111111111111110000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111000000000000001111111111111111111111111100000000000000000000000000011111111111110000000000000000000111100000000000000000001111111111111110000000000000000000000000001111111111111111111100000000000000000000000000001111111111111000000000000000000111100000000000000000000111111111111100000000000001111111111111110000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111100000000000111111111111111111111111111000000000000000000000000000111111111111110000000000000000000111100000000000000000001111111111111111000000000000000000000000000111111111111111111100000000000000000000000000011111111111111000000000000000000111100000000000000000000111111111111100000000000001111111110000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111000000111111111111111111000000000000000000000000000000000000001111111111111110000000000000000000111100000000000000000001111111111111111110000000000000000000000000001111111111111110000000000000000000000000000111111111111111000000000000000000111100000000000000000000111111111111100000000000001111000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000111100000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111110000000000000000000111100000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000111100000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000111111111111111111110000000000000000000111100000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000111100000000000000000000111111111111000000000000001111111111111111110000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111110000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111000000001111111111111111111111111111100000000000000000000000000000000111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000111111111111111111110000000000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000111111111111000011111111111111111111111111111111111000000000000000000000000000000011111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111110000000000000000000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111110000000000000000000000000000001111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000001111111111111110000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111110000000001111111111111111111111111110000000000000000000000000000011111111111110000000000000000000111100000000000000000001111111111111111100000000000000000000000000011111111111111110000000000000000000000000000011111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111000000000000001111111111111111111111111100000000000000000000000000001111111111110000000000000000000111100000000000000000001111111111111111000000000000000000000000001111111111111111111100000000000000000000000000001111111111111000000000000000000111100000000000000000000111111111111111111000000011111111111111111111111111111100000000000000000000000000000111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000011111111111111111111111110000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111100000000000000000000000000001111111111111111111100000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000001111111111111111111111110000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000011111111111111111111110000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111100000000000000000111111111111111111111111110000000000000000000000000000111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000111111111111111111111110000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000011111111111111111111110000000000000000000000000000011111111111000000000000000000111100000000000000000000111111111111000000000000000000011111111111111111111111100000000000000000000000000001111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111000000000000000000000001111111111111111111110000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000011111111111111111111110000000000000000000000000000011111111111000000000000000000111100000000000000000000111111111110000000000000000000001111111111111111111111100000000000000000000000000001111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000111111111111111111100000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000001111111111111111111100000000000000000000000000000011111111111000000000000000000111100000000000000000000111111111110000000000000000000000111111111111111111111000000000000000000000000000001111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000001111111111111110000000000000000000000000000000011111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000000111111111111111111000000000000000000000000000000011111111111000000000000000000111100000000000000000000111111111110000000000000000000000011111111111111111100000000000000000000000000000011111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111000000000000000000000000000000001111111111111100000000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111110000000000000000000000000111111111111100000000000000000000000000000000111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000111100000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000111100000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000111100000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000111100000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000111100000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000111100000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000111100000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000111100000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000111100000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000111100000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000011000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111100000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000111100000000000000000000111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000001100000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111110000000000000000000111100000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000111100000000000000000000111111111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000001111111111111111111111111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111110000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111100000000000000000000111100000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000111100000000000000000000011111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000001111111111111111111111111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000011000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000011000000000000000000000000111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000111111111111111111111111110000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000011111111111111111111111111111100000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000011111111111111111111111111111100000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001,
		512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
		512'b10010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001,
		512'b11010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001,
		512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
	 };
	 always_comb begin
		data[0]  = ROM[addr - 7];
		data[1]  = ROM[addr - 6];
		data[2]  = ROM[addr - 5];
		data[3]  = ROM[addr - 4];
		data[4]  = ROM[addr - 3];
		data[5]  = ROM[addr - 2];
		data[6]  = ROM[addr - 1];
		data[7]  = ROM[addr];
		data[8]  = ROM[addr + 1];
		data[9]  = ROM[addr + 2];
		data[10] = ROM[addr + 3];
		data[11] = ROM[addr + 4];
		data[12] = ROM[addr + 5];
		data[13] = ROM[addr + 6];
		data[14] = ROM[addr + 7];
		data[15] = ROM[addr + 8];
	 end
endmodule 