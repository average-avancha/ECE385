module mapROM  (input  [8:0] addr, 
                output [511:0] data);
    parameter ADDR_WIDTH = 9;
    parameter DATA_WIDTH = 512;
    
    parameter [0:2**ADDR_WIDTH - 1][DATA_WIDTH-1:0] ROM = {
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111110,
512'b01111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111,
512'b00111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111110,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111100000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000011111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111110,
512'b01111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111,
512'b01100000000000000000000000000000000000000000001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01111111111111111111111111111111111111111110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111,
512'b00111111111111111111111111111111111111111110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111110,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000011111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000001111110000000111111000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000011111110000000111111000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011100000000000000000000110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011110000000000000111100000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000111110000000000000111110000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011100000000000000000000110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000111000000000000000001110000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000001111000000000000000001110000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011100000000000000000000110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000001110000000000000000000111000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000001110000001111110000000111000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011100000000000000000001110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000011100000011111100000000111000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000011100000011111111100000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011000000000000000000001110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000011100000111111111000000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000011000000111000111110000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011000000111111111111111110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000111000001111000111100000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000001110000001110000001100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011000001111111111111111110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000111111111100000011100000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000001110000000110000001100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011000001100000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000111111111100000001100000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000001110000000111000001100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011000001100000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011111000000001110000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000110000001110000000111000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011000011100000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000001100000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000000111000000110000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000011100111111110000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000011100000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000000011110001110000011000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000011111111111111100000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000111100000111000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000000001111111110001111000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000001111110000011111000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000111111111000001111000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000011100000000011111100011110000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000000110000000000111100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000111111100000011110000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000011100000000000110000011100000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000000000000000000011110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000110000000000111100000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000001110000000000000000111000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000000000000000000001110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000110000000000110000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000111000000000000000011110000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000000011111100000000111000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000110000000000111100000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000011100000000000000001111000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111111001111111110000000011000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000110000000000011110000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000001111000000000000000000111000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111111111110001111000000011100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000111111110000000111000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000011110000011100000000000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000001111111000000011100000011100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000111111111000000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111100000111111100000000001110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000001100000001100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000011100000001110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000001110111111000000001110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000001100000001100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000001110000001110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001110000011100001111100000000110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000001110000001100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000001111111000000000110000001110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001110000011000000001110000000110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111111110000000001110000001100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000011111111111000000000110000000110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001100000011000000000110000000110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000011111111110000000001100000001100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000001111111011000000000110000000110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001100000011000000000111000000110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000011111110111000000001100000011100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000001110000011100000001110000001110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001100000011000000000111000000110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000001100000011100000011100000011100000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000001110000001111000111100000001110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001110000011100000000110000001110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000001110000011110001111000000011000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000111000000111111111000000001110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000001110000001111000011110000001110000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000001110000001111111110000000111000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000111000000011111110000000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000110000000111111111100000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000111000000011111100000001110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000011100000000000000000000011100000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000111000000001111111000000011100000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011100000000000000000001110000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000001111000000000000000001111000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000011100000000000000000001111000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011110000000000000000111100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000111100000000000000011110000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000001111000000000000000111110000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000001111100000000000001111000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011111110000000111111100000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000111111100000001111111100000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000011111100000011111110000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111110,
512'b01111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111,
512'b00111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111100000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000011111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111110,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111110,
512'b01111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01100000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000011,
512'b01111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111,
512'b00111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111110,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000110000000000000000110000000000000000000110000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111110000000000000000111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111100000000000000000011111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001100000000000000001100000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011000000000000000011000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    assign data = ROM[addr];
endmodule 